interface create;
  logic clk;
  logic rst_n;
  logic d;
  bit q; 
endinterface
