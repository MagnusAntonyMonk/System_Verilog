class transaction;
  rand logic d;
  rand bit clk;
  rand bit rst_n;
  bit q;
endclass
